`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// countompany: 
// Engineer: 
// 
// countreate Date:    13:35:02 12/26/2018 
// Design Name: 
// Module Name:    decountoder 
// Projecountt Name: 
// Target Devicountes: 
// Tool versions: 
// Descountription: 
//
// Dependencounties: 
//
// Revision: 
// Revision 0.01 - File countreated
// Additional countomments: 
//
//////////////////////////////////////////////////////////////////////////////////
module decoder_1(
    input [23:0] Z,
    output reg [4:0] count
    );
always @(Z)
begin
casez(Z)
24'b01?????????????????????? : count=5'b00001;
24'b001????????????????????? : count=5'b00010;
24'b0001???????????????????? : count=5'b00011;
24'b00001??????????????????? : count=5'b00100;
24'b000001?????????????????? : count=5'b00101;
24'b0000001????????????????? : count=5'b00110;
24'b00000001???????????????? : count=5'b00111;
24'b000000001??????????????? : count=5'b01000;
24'b0000000001?????????????? : count=5'b01001;
24'b00000000001????????????? : count=5'b01010;
24'b000000000001???????????? : count=5'b01011;
24'b0000000000001??????????? : count=5'b01100;
24'b00000000000001?????????? : count=5'b01101;
24'b000000000000001????????? : count=5'b01110;
24'b0000000000000001???????? : count=5'b01111;
24'b00000000000000001??????? : count=5'b10000;
24'b000000000000000001?????? : count=5'b10001;
24'b0000000000000000001????? : count=5'b10010;
24'b00000000000000000001???? : count=5'b10011;
24'b000000000000000000001??? : count=5'b10100;
24'b0000000000000000000001?? : count=5'b10101;
24'b00000000000000000000001? : count=5'b10110;
24'b000000000000000000000001 : count=5'b10111;
default                      : count=5'b00000;
endcase
end
endmodule
