`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:49:14 08/07/2019 
// Design Name: 
// Module Name:    adder12 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module adder9(
    input [8:0] a,
    input [8:0] b,
    output [8:0] s
    );

assign s=a+b;

endmodule
