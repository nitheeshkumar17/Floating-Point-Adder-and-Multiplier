`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:48:14 08/07/2019 
// Design Name: 
// Module Name:    adder6 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module adder6(
    input [5:0] a,
    input [5:0] b,
    output [5:0] s
    );

assign s=a+b;

endmodule
